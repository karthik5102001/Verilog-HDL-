module Testing_iverilog (A,b);
input A;
output b;

assign b =~ A;

endmodule